magic
tech scmos
timestamp 1481247542
<< nwell >>
rect -25 -17 27 41
<< ptransistor >>
rect -8 -9 -6 23
rect 0 -9 2 23
rect 8 -9 10 23
<< pdiffusion >>
rect -9 -9 -8 23
rect -6 -9 -5 23
rect -1 -9 0 23
rect 2 -9 3 23
rect 7 -9 8 23
rect 10 -9 11 23
<< pdcontact >>
rect -13 -9 -9 23
rect -5 -9 -1 23
rect 3 -9 7 23
rect 11 -9 15 23
<< nsubstratencontact >>
rect -19 34 21 38
<< polysilicon >>
rect -8 24 10 26
rect -8 23 -6 24
rect 0 23 2 24
rect 8 23 10 24
rect -8 -11 -6 -9
rect 0 -11 2 -9
rect 8 -11 10 -9
<< polycontact >>
rect -1 26 3 30
<< metal1 >>
rect -23 38 25 39
rect -23 34 -19 38
rect 21 34 25 38
rect -23 33 25 34
rect -13 23 -9 33
rect 11 23 15 33
rect -5 -12 -1 -9
rect -15 -16 -1 -12
rect 3 -12 7 -9
rect 3 -16 17 -12
<< m2contact >>
rect 3 26 7 30
rect -19 -16 -15 -12
rect 17 -16 21 -12
<< metal2 >>
rect -19 -20 -15 -16
rect 17 -20 21 -16
<< labels >>
rlabel m2contact 5 28 5 28 1 Clk
rlabel metal2 -17 -18 -17 -18 1 Bl
rlabel metal2 19 -18 19 -18 1 Bl_
<< end >>
