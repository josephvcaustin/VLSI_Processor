magic
tech scmos
timestamp 1481316610
<< error_s >>
rect 227 452 233 454
<< nwell >>
rect 904 1174 927 1178
<< metal1 >>
rect -168 1237 1095 1252
rect -168 451 -153 1237
rect 514 1166 532 1237
rect 944 1172 958 1237
rect 1080 492 1095 1237
rect 958 478 1095 492
rect -168 436 266 451
rect -168 218 -153 436
rect 597 327 601 378
rect 644 334 648 378
rect 691 341 695 378
rect 738 348 742 378
rect 785 355 789 378
rect 832 362 836 378
rect 879 369 883 378
rect 926 376 930 379
rect 926 372 1042 376
rect 879 365 1035 369
rect 832 358 1028 362
rect 785 351 1021 355
rect 738 344 1014 348
rect 691 337 1007 341
rect 644 330 1000 334
rect 597 323 993 327
rect -168 200 -19 218
rect -168 -338 -153 200
rect 989 108 993 323
rect 662 104 993 108
rect 662 62 666 104
rect 996 101 1000 330
rect 710 97 1000 101
rect 710 61 714 97
rect 1003 94 1007 337
rect 758 90 1007 94
rect 758 61 762 90
rect 1010 87 1014 344
rect 814 83 1014 87
rect 1017 80 1021 351
rect 861 76 1021 80
rect 1024 73 1028 358
rect 908 69 1028 73
rect 1031 66 1035 365
rect 955 62 1035 66
rect 1038 59 1042 372
rect 1002 55 1042 59
rect 637 45 642 52
rect 1080 -39 1095 478
rect 617 -40 660 -39
rect 617 -43 664 -40
rect 1021 -43 1095 -39
rect 617 -46 660 -43
rect 1022 -46 1095 -43
rect 617 -96 624 -46
rect 1080 -96 1095 -46
rect 617 -103 644 -96
rect 1022 -103 1095 -96
rect 617 -195 624 -103
rect 639 -146 643 -139
rect 1080 -195 1095 -103
rect 617 -198 642 -195
rect 617 -200 651 -198
rect 617 -204 639 -200
rect 643 -204 651 -200
rect 617 -205 651 -204
rect 1022 -205 1095 -195
rect 617 -208 642 -205
rect 1022 -206 1025 -205
rect 617 -315 624 -208
rect 1021 -209 1025 -206
rect 1029 -209 1095 -205
rect 637 -263 642 -256
rect 617 -321 643 -315
rect 1014 -321 1018 -319
rect 617 -338 624 -321
rect 1014 -338 1022 -321
rect 1080 -338 1095 -209
rect -168 -353 1095 -338
<< m2contact >>
rect 923 1174 927 1178
rect 597 378 601 382
rect 644 378 648 382
rect 691 378 695 382
rect 738 378 742 382
rect 785 378 789 382
rect 832 378 836 382
rect 879 378 883 382
rect 926 379 930 383
rect 11 313 15 317
rect 136 313 140 317
rect 261 313 265 317
rect 386 313 390 317
rect 511 313 515 317
rect 636 313 640 317
rect 761 313 765 317
rect 886 314 890 318
rect -20 306 -13 313
rect 982 156 986 160
rect -23 111 -15 119
rect 662 58 666 62
rect 710 57 714 61
rect 810 83 814 87
rect 857 76 861 80
rect 904 69 908 73
rect 951 62 955 66
rect 758 57 762 61
rect 998 55 1002 59
rect 631 45 637 52
rect 1021 45 1027 52
rect 633 -146 639 -139
rect 1021 -146 1027 -139
rect 639 -204 643 -200
rect 1025 -209 1029 -205
rect 631 -263 637 -256
rect 1021 -263 1027 -256
<< metal2 >>
rect 1105 1277 1120 1278
rect -194 1262 1120 1277
rect -193 452 -178 1262
rect 198 1203 210 1262
rect 532 1189 547 1262
rect 904 1174 923 1178
rect 959 1154 971 1262
rect 1105 590 1120 1262
rect 971 578 1120 590
rect -193 440 200 452
rect -193 313 -178 440
rect -16 386 31 390
rect -16 377 24 381
rect -16 368 17 372
rect -16 358 10 362
rect 6 353 10 358
rect 13 360 17 368
rect 20 367 24 377
rect 27 374 31 386
rect 27 370 878 374
rect 20 363 753 367
rect 13 356 628 360
rect -16 349 3 353
rect 6 349 503 353
rect -1 346 3 349
rect -16 340 -4 344
rect -1 342 378 346
rect -8 339 -4 340
rect -8 335 253 339
rect -16 332 -11 334
rect -16 330 128 332
rect -15 328 128 330
rect -16 324 3 325
rect -16 321 -1 324
rect 124 324 128 328
rect 249 321 253 335
rect 374 317 378 342
rect 499 318 503 349
rect 624 313 628 356
rect 749 315 753 363
rect 874 324 878 370
rect -193 306 -20 313
rect -193 119 -178 306
rect 974 150 978 156
rect -10 137 -3 141
rect -193 111 -23 119
rect -193 -363 -178 111
rect -7 86 -3 137
rect 849 111 853 113
rect 849 109 932 111
rect 853 107 932 109
rect 99 69 103 107
rect 224 76 228 107
rect 349 83 353 107
rect 474 90 478 107
rect 599 97 603 107
rect 724 104 728 107
rect 724 100 885 104
rect 599 93 837 97
rect 474 86 790 90
rect 349 79 742 83
rect 224 72 694 76
rect 99 65 646 69
rect 642 57 646 65
rect 624 52 635 54
rect 690 57 694 72
rect 738 57 742 79
rect 786 57 790 86
rect 833 57 837 93
rect 880 57 884 100
rect 927 57 931 107
rect 974 57 978 114
rect 1105 52 1120 578
rect 624 45 631 52
rect 1027 45 1120 52
rect 624 -139 635 45
rect 679 36 1013 40
rect 1105 -139 1120 45
rect 624 -146 633 -139
rect 1027 -146 1120 -139
rect 624 -256 635 -146
rect 1105 -256 1120 -146
rect 624 -263 631 -256
rect 1027 -263 1120 -256
rect 624 -363 635 -263
rect 660 -312 1064 -308
rect 1105 -363 1120 -263
rect -193 -378 1120 -363
<< m3contact >>
rect 927 1174 931 1178
rect 950 399 954 403
rect -20 386 -16 390
rect -20 377 -16 381
rect -20 368 -16 372
rect -20 358 -16 362
rect 597 382 601 386
rect 644 382 648 386
rect 691 382 695 386
rect 738 382 742 386
rect 785 382 789 386
rect 832 382 836 386
rect 879 382 883 386
rect 926 383 930 387
rect -20 349 -16 353
rect -20 340 -16 344
rect -20 330 -16 334
rect -20 321 -16 325
rect 31 321 35 325
rect 156 321 160 325
rect 281 321 285 325
rect 406 321 410 325
rect 531 321 535 325
rect 656 321 660 325
rect 781 322 785 326
rect 906 320 910 324
rect 986 156 990 160
rect 642 53 646 57
rect 662 54 666 58
rect 690 53 694 57
rect 710 53 714 57
rect 738 53 742 57
rect 758 53 762 57
rect 806 83 810 87
rect 786 53 790 57
rect 853 76 857 80
rect 833 53 837 57
rect 900 69 904 73
rect 880 53 884 57
rect 947 62 951 66
rect 927 53 931 57
rect 974 53 978 57
rect 994 53 998 59
rect 639 -208 643 -204
rect 1021 -209 1025 -205
rect 1064 -312 1068 -308
<< metal3 >>
rect -199 1186 190 1192
rect 926 1178 1126 1179
rect -199 1172 189 1178
rect 926 1174 927 1178
rect 931 1174 1126 1178
rect 926 1173 1126 1174
rect -199 1156 190 1162
rect 498 1101 504 1107
rect 498 1057 504 1063
rect 498 951 504 957
rect 498 891 504 897
rect -199 815 192 821
rect -199 801 190 807
rect 498 801 504 807
rect -199 785 190 791
rect 498 711 504 717
rect 498 621 504 627
rect 964 567 1126 573
rect 498 528 504 534
rect 949 403 1126 404
rect 949 399 950 403
rect 954 399 1126 403
rect 949 398 1126 399
rect -199 390 -15 391
rect -199 386 -20 390
rect -16 386 -15 390
rect -199 385 -15 386
rect -199 381 -15 382
rect 576 381 582 387
rect -199 377 -20 381
rect -16 377 -15 381
rect -199 376 -15 377
rect 30 375 582 381
rect -199 372 -15 373
rect -199 368 -20 372
rect -16 368 -15 372
rect -199 367 -15 368
rect -199 362 -15 363
rect -199 358 -20 362
rect -16 358 -15 362
rect -199 357 -15 358
rect -199 353 -15 354
rect -199 349 -20 353
rect -16 349 -15 353
rect -199 348 -15 349
rect -199 344 -15 345
rect -199 340 -20 344
rect -16 340 -15 344
rect -199 339 -15 340
rect -199 334 -15 335
rect -199 330 -20 334
rect -16 330 -15 334
rect -199 329 -15 330
rect -199 325 -15 326
rect -199 321 -20 325
rect -16 321 -15 325
rect -199 320 -15 321
rect 30 325 36 375
rect 623 372 629 386
rect 30 321 31 325
rect 35 321 36 325
rect 30 320 36 321
rect 155 366 629 372
rect 155 325 161 366
rect 670 363 676 387
rect 155 321 156 325
rect 160 321 161 325
rect 155 320 161 321
rect 280 357 676 363
rect 280 325 286 357
rect 717 354 723 387
rect 280 321 281 325
rect 285 321 286 325
rect 280 320 286 321
rect 405 348 723 354
rect 405 325 411 348
rect 764 345 770 387
rect 405 321 406 325
rect 410 321 411 325
rect 405 320 411 321
rect 530 339 770 345
rect 530 325 536 339
rect 811 336 817 387
rect 530 321 531 325
rect 535 321 536 325
rect 530 320 536 321
rect 655 330 817 336
rect 655 325 661 330
rect 858 327 864 387
rect 655 321 656 325
rect 660 321 661 325
rect 780 326 864 327
rect 780 322 781 326
rect 785 322 864 326
rect 780 321 864 322
rect 905 324 911 388
rect 655 320 661 321
rect 905 320 906 324
rect 910 320 911 324
rect 905 319 911 320
rect -199 273 -17 279
rect 985 273 1000 279
rect -199 253 -19 259
rect 994 161 1000 273
rect 982 160 1000 161
rect 982 156 986 160
rect 990 156 1000 160
rect 982 155 1000 156
rect 805 87 811 88
rect 805 83 806 87
rect 810 83 811 87
rect 661 58 667 59
rect 641 57 647 58
rect 641 53 642 57
rect 646 53 647 57
rect 641 -125 647 53
rect 661 54 662 58
rect 666 54 667 58
rect 661 2 667 54
rect 689 57 695 58
rect 689 53 690 57
rect 694 53 695 57
rect 689 -125 695 53
rect 709 57 715 58
rect 709 53 710 57
rect 714 53 715 57
rect 709 2 715 53
rect 737 57 743 58
rect 737 53 738 57
rect 742 53 743 57
rect 737 -125 743 53
rect 757 57 763 58
rect 757 53 758 57
rect 762 53 763 57
rect 757 2 763 53
rect 785 57 791 58
rect 785 53 786 57
rect 790 53 791 57
rect 785 -125 791 53
rect 805 2 811 83
rect 852 80 858 81
rect 852 76 853 80
rect 857 76 858 80
rect 832 57 838 58
rect 832 53 833 57
rect 837 53 838 57
rect 832 -125 838 53
rect 852 2 858 76
rect 899 73 905 74
rect 899 69 900 73
rect 904 69 905 73
rect 879 57 885 58
rect 879 53 880 57
rect 884 53 885 57
rect 879 -125 885 53
rect 899 2 905 69
rect 946 66 952 67
rect 946 62 947 66
rect 951 62 952 66
rect 926 57 932 58
rect 926 53 927 57
rect 931 53 932 57
rect 926 -125 932 53
rect 946 2 952 62
rect 993 59 999 60
rect 973 57 979 58
rect 973 53 974 57
rect 978 53 979 57
rect 973 -125 979 53
rect 993 53 994 59
rect 998 53 999 59
rect 993 2 999 53
rect 1011 35 1126 41
rect 1017 -134 1126 -128
rect 638 -204 648 -203
rect 638 -208 639 -204
rect 643 -208 648 -204
rect 638 -209 648 -208
rect 642 -258 648 -209
rect 1016 -205 1026 -204
rect 1016 -209 1021 -205
rect 1025 -209 1026 -205
rect 1016 -210 1026 -209
rect 1016 -252 1022 -210
rect 1017 -257 1022 -252
rect 1063 -308 1126 -307
rect 1063 -312 1064 -308
rect 1068 -312 1126 -308
rect 1063 -313 1126 -312
use rf_dec  rf_dec_0
timestamp 1481316610
transform 1 0 553 0 1 399
box -364 -19 418 811
use alu  alu_0
timestamp 1481316610
transform 1 0 -21 0 1 51
box 1 56 1007 273
use alu_reg  alu_reg_0
timestamp 1481316610
transform -1 0 1021 0 -1 15
box -4 -37 381 338
<< labels >>
rlabel metal3 -199 253 -193 259 7 Select
rlabel metal3 -199 273 -193 279 7 Subtract
rlabel metal3 -199 320 -193 326 7 I7
rlabel metal3 -199 329 -193 335 7 I6
rlabel metal3 -199 339 -193 345 7 I5
rlabel metal3 -199 348 -193 354 7 I4
rlabel metal3 -199 357 -193 363 7 I3
rlabel metal3 -199 367 -193 373 7 I2
rlabel metal3 -199 376 -193 382 7 I1
rlabel metal3 -199 385 -193 391 7 I0
rlabel metal3 1120 -134 1126 -128 7 ALU_Ds
rlabel metal3 1120 35 1126 41 7 ALU_As
rlabel metal3 1120 398 1126 404 3 REG_As
rlabel metal3 1120 567 1126 573 3 REG_Ds
rlabel metal3 1120 1173 1126 1179 3 REG_Pc
rlabel metal3 -199 1156 -193 1162 7 A0
rlabel metal3 -199 1172 -193 1178 7 A1
rlabel metal3 -199 1186 -193 1192 7 A2
rlabel metal3 -199 785 -193 791 7 D0
rlabel metal3 -199 801 -193 807 7 D1
rlabel metal3 -199 815 -193 821 7 D2
rlabel metal3 1120 -313 1126 -307 3 ALU_Pc
rlabel metal1 989 108 993 112 1 O7
rlabel metal1 996 108 1000 112 1 O6
rlabel metal1 1003 108 1007 112 1 O5
rlabel metal1 1010 108 1014 112 1 O4
rlabel metal1 1017 108 1021 112 1 O3
rlabel metal1 1024 108 1028 112 1 O2
rlabel metal1 1031 108 1035 112 1 O1
rlabel metal1 1038 108 1042 112 1 O0
rlabel metal2 458 1262 498 1277 0 gnd
rlabel metal1 458 1237 498 1252 0 vdd
rlabel metal3 576 381 582 387 5 Ad7
rlabel metal3 623 380 629 386 5 Ad6
rlabel metal3 670 381 676 387 5 Ad5
rlabel metal3 717 381 723 387 5 Ad4
rlabel metal3 764 381 770 387 5 Ad3
rlabel metal3 811 381 817 387 5 Ad2
rlabel metal3 858 381 864 387 5 Ad1
rlabel metal3 905 382 911 388 5 Ad0
rlabel metal2 99 91 103 95 1 S7
rlabel metal2 224 93 228 97 1 S6
rlabel metal2 349 93 353 97 1 S5
rlabel metal2 474 96 478 100 1 S4
rlabel metal2 599 99 603 103 1 S3
rlabel metal2 724 101 728 104 1 S2
rlabel metal2 856 108 860 111 1 S1
rlabel metal2 974 108 978 111 1 S0
rlabel metal2 -7 86 -3 90 1 S8
rlabel metal3 498 1101 504 1107 1 En0
rlabel metal3 498 1057 504 1063 1 En1
rlabel metal3 498 951 504 957 1 En2
rlabel metal3 498 891 504 897 1 En3
rlabel metal3 498 801 504 807 1 En4
rlabel metal3 498 711 504 717 1 En5
rlabel metal3 498 621 504 627 1 En6
rlabel metal3 498 528 504 534 1 En7
<< end >>
