magic
tech scmos
timestamp 1480717170
<< ntransistor >>
rect -3 -55 -1 -25
rect 5 -55 7 -25
rect 21 -55 23 -45
<< ptransistor >>
rect -3 0 -1 30
rect 5 0 7 30
rect 21 10 23 30
<< ndiffusion >>
rect -4 -55 -3 -25
rect -1 -55 0 -25
rect 4 -55 5 -25
rect 7 -55 8 -25
rect 20 -55 21 -45
rect 23 -55 24 -45
<< pdiffusion >>
rect -4 0 -3 30
rect -1 0 0 30
rect 4 0 5 30
rect 7 0 8 30
rect 20 10 21 30
rect 23 10 24 30
<< ndcontact >>
rect -8 -55 -4 -25
rect 0 -55 4 -25
rect 8 -55 12 -25
rect 16 -55 20 -45
rect 24 -55 28 -45
<< pdcontact >>
rect -8 0 -4 30
rect 0 0 4 30
rect 8 0 12 30
rect 16 10 20 30
rect 24 10 28 30
<< psubstratepcontact >>
rect -8 -68 28 -62
<< nsubstratencontact >>
rect -8 34 28 40
<< polysilicon >>
rect -3 30 -1 32
rect 5 30 7 32
rect 21 30 23 32
rect -3 -7 -1 0
rect 5 -14 7 0
rect 21 -7 23 10
rect -3 -17 4 -15
rect -3 -25 -1 -17
rect 21 -22 23 -11
rect 5 -24 23 -22
rect 5 -25 7 -24
rect 21 -45 23 -24
rect -3 -57 -1 -55
rect 5 -57 7 -55
rect 21 -57 23 -55
<< polycontact >>
rect -4 -11 0 -7
rect 20 -11 24 -7
rect 4 -18 8 -14
<< metal1 >>
rect -12 40 32 41
rect -12 34 -8 40
rect 28 34 32 40
rect -12 33 32 34
rect 24 30 28 33
rect 0 -11 20 -7
rect 8 -18 16 -14
rect 16 -45 20 -18
rect 24 -62 28 -55
rect -12 -68 -8 -62
rect 28 -68 32 -62
rect -12 -69 32 -68
<< m2contact >>
rect -8 -4 -4 0
rect 0 -4 4 0
rect 16 6 20 10
rect 8 -4 12 0
rect 16 -18 20 -14
rect -8 -25 -4 -21
rect 0 -25 4 -21
rect 8 -25 12 -21
<< metal2 >>
rect -8 -21 -4 -4
rect 0 -21 4 -4
rect 8 -21 12 -4
rect 16 -14 20 6
<< labels >>
rlabel psubstratepcontact 10 -65 10 -65 0 GND
rlabel nsubstratencontact 10 37 10 37 0 VDD
rlabel metal1 14 -9 14 -9 0 S
rlabel metal2 10 -13 10 -13 0 B
rlabel metal2 -6 -14 -6 -14 0 A
rlabel metal2 2 -13 2 -13 0 OUT
<< end >>
