magic
tech scmos
timestamp 1480732973
<< nwell >>
rect -13 -10 38 16
<< ntransistor >>
rect 5 -25 7 -17
rect 21 -25 23 -17
rect -2 -32 4 -30
rect 24 -32 30 -30
<< ptransistor >>
rect 5 0 7 4
rect 21 0 23 4
<< ndiffusion >>
rect 4 -25 5 -17
rect 7 -25 8 -17
rect 20 -25 21 -17
rect 23 -25 24 -17
rect -2 -30 4 -28
rect -2 -33 4 -32
rect 24 -30 30 -28
rect 24 -33 30 -32
<< pdiffusion >>
rect 4 0 5 4
rect 7 0 8 4
rect 20 0 21 4
rect 23 0 24 4
<< ndcontact >>
rect -2 -28 4 -17
rect 8 -25 12 -17
rect 16 -25 20 -17
rect 24 -28 30 -17
rect -2 -37 4 -33
rect 24 -37 30 -33
<< pdcontact >>
rect 0 0 4 4
rect 8 0 12 4
rect 16 0 20 4
rect 24 0 28 4
<< psubstratepcontact >>
rect -6 -45 3 -41
rect 13 -45 34 -41
<< nsubstratencontact >>
rect -6 8 34 12
<< polysilicon >>
rect 5 4 7 6
rect 21 4 23 6
rect 5 -17 7 0
rect 21 -17 23 0
rect 5 -27 7 -25
rect 21 -27 23 -25
rect -4 -32 -2 -30
rect 4 -32 13 -30
rect 17 -32 24 -30
rect 30 -32 32 -30
<< polycontact >>
rect 17 -7 21 -3
rect 7 -14 11 -10
rect 13 -33 17 -29
<< metal1 >>
rect -10 12 38 14
rect -10 8 -6 12
rect 34 8 38 12
rect -10 7 38 8
rect 8 4 12 7
rect 16 4 20 7
rect 0 -3 4 0
rect 0 -7 17 -3
rect 0 -17 4 -7
rect 24 -10 28 0
rect 11 -14 28 -10
rect 24 -17 28 -14
rect 13 -37 17 -33
rect -10 -41 6 -40
rect -10 -45 -6 -41
rect 3 -45 6 -41
rect 10 -41 38 -40
rect 10 -45 13 -41
rect 34 -45 38 -41
rect -10 -47 38 -45
<< m2contact >>
rect 12 -25 16 -17
rect -6 -37 -2 -33
rect 17 -37 21 -33
rect 30 -37 34 -33
rect 6 -45 10 -40
<< metal2 >>
rect -6 -33 -2 14
rect -6 -47 -2 -37
rect 6 -25 12 -17
rect 6 -40 10 -25
rect 30 -33 34 14
rect 30 -47 34 -37
<< m3contact >>
rect 17 -41 21 -37
<< metal3 >>
rect -10 -37 38 -36
rect -10 -41 17 -37
rect 21 -41 38 -37
rect -10 -42 38 -41
<< labels >>
rlabel nsubstratencontact 14 10 14 10 1 Vdd
rlabel metal1 12 -44 12 -44 1 Gnd
rlabel metal3 36 -39 36 -39 1 En
rlabel metal2 -4 -23 -4 -23 1 Bl
rlabel metal2 32 -23 32 -23 1 Bl_
<< end >>
