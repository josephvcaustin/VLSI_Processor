magic
tech scmos
timestamp 1481248605
<< nwell >>
rect 43 782 51 788
rect 4 733 8 737
rect 333 733 337 737
rect 163 36 173 38
<< metal1 >>
rect -155 805 -149 806
rect -277 799 -21 805
rect -277 781 -271 799
rect -220 787 -214 789
rect -39 730 -21 799
rect 396 788 405 799
rect 43 782 51 788
rect 392 782 405 788
rect 391 730 405 782
rect -39 723 1 730
rect 374 723 405 730
rect -39 699 -21 723
rect -51 692 -21 699
rect -59 688 -21 692
rect -51 681 -21 688
rect -39 615 -21 681
rect 376 615 381 616
rect 391 615 405 723
rect -39 601 1 615
rect 376 601 405 615
rect -39 519 -21 601
rect -55 501 -21 519
rect -39 493 -21 501
rect 391 493 405 601
rect -39 479 2 493
rect 377 479 405 493
rect -39 371 -21 479
rect 391 371 405 479
rect -39 357 1 371
rect 376 357 405 371
rect -39 339 -21 357
rect -52 321 -21 339
rect -39 249 -21 321
rect 391 249 405 357
rect -39 235 0 249
rect 377 235 405 249
rect -39 159 -21 235
rect -51 143 -21 159
rect 391 143 405 235
rect -51 141 0 143
rect -39 136 0 141
rect 376 136 405 143
rect -287 52 -272 75
rect -221 69 -215 115
rect -39 86 -21 136
rect 391 86 405 136
rect -39 79 1 86
rect 376 85 405 86
rect 375 79 405 85
rect -221 60 -135 69
rect -39 52 -21 79
rect -287 37 -21 52
rect -39 -13 -21 37
<< m2contact >>
rect -220 789 -214 794
rect -51 771 -45 780
rect 4 733 8 737
rect 333 733 337 737
rect -58 703 -54 707
rect -58 659 -54 663
rect -6 662 0 676
rect 377 662 384 676
rect -53 591 -47 609
rect -59 553 -55 557
rect -6 539 0 554
rect 377 540 384 554
rect -58 493 -54 497
rect -331 431 -325 443
rect -51 411 -45 429
rect -58 403 -54 407
rect -6 419 0 432
rect 377 418 384 432
rect -58 313 -54 317
rect -7 296 0 310
rect 377 296 384 310
rect -55 231 -48 249
rect -58 223 -54 227
rect -7 179 0 186
rect 376 179 383 186
rect -58 130 -54 134
rect -326 53 -320 60
rect -55 61 -48 68
rect -3 -12 4 -5
<< metal2 >>
rect -355 443 -343 811
rect -21 794 -6 796
rect -214 789 -6 794
rect 411 792 418 799
rect -21 780 -6 789
rect -45 771 -6 780
rect 22 775 26 779
rect -50 770 -6 771
rect -21 680 -6 770
rect -21 676 -3 680
rect 406 676 418 792
rect -21 609 -6 676
rect 384 662 418 676
rect -47 591 -6 609
rect -355 431 -331 443
rect -355 53 -343 431
rect -21 429 -6 591
rect 406 554 418 662
rect 384 540 418 554
rect 406 432 418 540
rect -45 411 -6 429
rect 384 418 418 432
rect -21 310 -6 411
rect 406 310 418 418
rect -21 296 -7 310
rect 384 296 418 310
rect -21 249 -6 296
rect -48 231 -6 249
rect -21 186 -6 231
rect 406 186 418 296
rect -21 179 -7 186
rect 383 179 418 186
rect -21 68 -6 179
rect -48 61 -6 68
rect -55 60 -6 61
rect -21 53 -6 60
rect -355 41 -6 53
rect -21 -5 -6 41
rect 0 0 401 4
rect -21 -12 -3 -5
rect -21 -13 4 -12
<< m3contact >>
rect -298 788 -294 792
rect -312 768 -308 772
rect -326 758 -322 762
rect -54 703 -50 707
rect -54 659 -50 663
rect -55 553 -51 557
rect -54 493 -50 497
rect -299 417 -295 421
rect -54 403 -50 407
rect -313 397 -309 401
rect -327 387 -323 391
rect -54 313 -50 317
rect -54 223 -50 227
rect -54 130 -50 134
<< metal3 >>
rect -363 792 -293 793
rect -363 788 -298 792
rect -294 788 -293 792
rect -363 787 -293 788
rect -152 781 -146 811
rect -142 781 -136 811
rect -364 773 -307 779
rect -315 772 -307 773
rect -315 768 -312 772
rect -308 768 -307 772
rect -315 767 -307 768
rect -364 762 -321 763
rect -364 758 -326 762
rect -322 758 -321 762
rect -364 757 -321 758
rect -55 707 -49 708
rect -55 703 -54 707
rect -50 703 -49 707
rect -55 680 -49 703
rect -55 674 6 680
rect -55 663 6 664
rect -55 659 -54 663
rect -50 659 6 663
rect -55 658 6 659
rect -56 557 6 558
rect -56 553 -55 557
rect -51 553 6 557
rect -56 552 6 553
rect -9 536 6 542
rect -9 498 -3 536
rect -55 497 -3 498
rect -55 493 -54 497
rect -50 493 -3 497
rect -55 492 -3 493
rect -9 491 -3 492
rect -38 430 6 436
rect -363 421 -294 422
rect -363 417 -299 421
rect -295 417 -294 421
rect -363 416 -294 417
rect -38 408 -32 430
rect -363 402 -308 408
rect -55 407 -32 408
rect -55 403 -54 407
rect -50 403 -32 407
rect -55 402 -32 403
rect -29 414 6 420
rect -314 401 -308 402
rect -314 397 -313 401
rect -309 397 -308 401
rect -314 396 -308 397
rect -363 391 -322 392
rect -363 387 -327 391
rect -323 387 -322 391
rect -363 386 -322 387
rect -29 318 -23 414
rect -55 317 -23 318
rect -55 313 -54 317
rect -50 313 -23 317
rect -55 312 -23 313
rect -20 308 6 314
rect -20 228 -14 308
rect -55 227 -14 228
rect -55 223 -54 227
rect -50 223 -14 227
rect -55 222 -14 223
rect -20 221 -14 222
rect -11 292 6 298
rect -11 135 -5 292
rect -55 134 -5 135
rect -55 130 -54 134
rect -50 130 -5 134
rect -55 129 -5 130
rect -1 75 5 174
rect 371 168 412 174
rect -152 9 -146 75
rect -143 69 5 75
rect -152 3 19 9
rect -152 2 -146 3
rect 23 -18 29 38
rect 43 -18 49 165
rect 70 -19 76 38
rect 90 -18 96 165
rect 117 -18 123 38
rect 137 -18 143 165
rect 164 -18 170 38
rect 184 -18 190 165
rect 211 -18 217 38
rect 231 -18 237 165
rect 258 -18 264 38
rect 278 -18 284 165
rect 305 -18 311 38
rect 325 -18 331 165
rect 342 127 348 134
rect 339 3 345 9
rect 352 -17 358 38
rect 372 -17 378 165
use decoder_full  decoder_full_0
timestamp 1481248605
transform 0 -1 -180 1 0 58
box -3 -129 731 147
use register_file  register_file_0
timestamp 1481247610
transform 1 0 -17 0 1 25
box 14 -37 396 765
<< labels >>
rlabel metal3 406 168 412 174 1 Ds
rlabel metal3 352 -17 358 -11 5 Ad0
rlabel metal3 372 -17 378 -11 5 Dd0
rlabel metal3 325 -18 331 -12 5 Dd1
rlabel metal3 305 -18 311 -12 5 Ad1
rlabel metal3 278 -18 284 -12 5 Dd2
rlabel metal3 258 -18 264 -12 5 Ad2
rlabel metal3 231 -18 237 -12 5 Dd3
rlabel metal3 211 -18 217 -12 5 Ad3
rlabel metal3 184 -18 190 -12 5 Dd4
rlabel metal3 164 -18 170 -12 5 Ad4
rlabel metal3 137 -18 143 -12 5 Dd5
rlabel metal3 117 -18 123 -12 5 Ad5
rlabel metal3 90 -18 96 -12 5 Dd6
rlabel metal3 70 -19 76 -13 5 Ad6
rlabel metal3 43 -18 49 -12 5 Dd7
rlabel metal3 23 -18 29 -12 5 Ad7
rlabel metal2 396 0 401 4 1 As
rlabel metal3 -364 757 -358 763 5 A0
rlabel metal3 -364 773 -358 779 5 A1
rlabel metal3 -363 787 -357 793 5 A2
rlabel metal3 -363 386 -357 392 5 D0
rlabel metal3 -363 402 -357 408 5 D1
rlabel metal3 -363 416 -357 422 5 D2
rlabel metal1 -28 799 -21 805 1 VDD
rlabel metal2 -13 790 -6 796 1 GND
rlabel metal3 -142 805 -136 811 1 Ds
rlabel metal3 -152 805 -146 811 1 As
rlabel metal3 342 128 348 134 5 iso_sel1
rlabel m2contact 333 733 337 737 1 Bl
rlabel metal1 45 782 50 788 1 PreV
rlabel metal2 22 775 26 779 1 Pc
<< end >>
