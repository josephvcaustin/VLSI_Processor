magic
tech scmos
timestamp 1480714837
<< ntransistor >>
rect -12 19 -10 29
rect -4 19 -2 29
rect 1 19 3 29
rect 9 19 11 29
rect 17 19 19 29
rect 25 19 27 29
rect 41 19 43 29
rect 49 19 51 29
rect 57 19 59 29
rect 65 19 67 29
rect 79 19 81 29
rect 84 19 86 29
rect 89 19 91 29
rect 97 19 99 29
<< ptransistor >>
rect -12 72 -10 92
rect -4 72 -2 92
rect 1 72 3 92
rect 9 72 11 92
rect 17 72 19 92
rect 25 72 27 92
rect 41 72 43 92
rect 49 72 51 92
rect 57 72 59 92
rect 65 72 67 92
rect 79 72 81 92
rect 84 72 86 92
rect 89 72 91 92
rect 97 72 99 92
<< ndiffusion >>
rect -13 19 -12 29
rect -10 19 -9 29
rect -5 19 -4 29
rect -2 19 1 29
rect 3 19 4 29
rect 8 19 9 29
rect 11 19 12 29
rect 16 19 17 29
rect 19 19 20 29
rect 24 19 25 29
rect 27 19 28 29
rect 40 19 41 29
rect 43 19 44 29
rect 48 19 49 29
rect 51 19 52 29
rect 56 19 57 29
rect 59 19 60 29
rect 64 19 65 29
rect 67 19 68 29
rect 78 19 79 29
rect 81 19 84 29
rect 86 19 89 29
rect 91 19 92 29
rect 96 19 97 29
rect 99 19 100 29
<< pdiffusion >>
rect -13 72 -12 92
rect -10 72 -9 92
rect -5 72 -4 92
rect -2 72 1 92
rect 3 72 4 92
rect 8 72 9 92
rect 11 72 12 92
rect 16 72 17 92
rect 19 72 20 92
rect 24 72 25 92
rect 27 72 28 92
rect 40 72 41 92
rect 43 72 44 92
rect 48 72 49 92
rect 51 72 52 92
rect 56 72 57 92
rect 59 72 60 92
rect 64 72 65 92
rect 67 72 68 92
rect 78 72 79 92
rect 81 72 84 92
rect 86 72 89 92
rect 91 72 92 92
rect 96 72 97 92
rect 99 72 100 92
<< ndcontact >>
rect -17 19 -13 29
rect -9 19 -5 29
rect 4 19 8 29
rect 12 19 16 29
rect 20 19 24 29
rect 28 19 32 29
rect 36 19 40 29
rect 44 19 48 29
rect 52 19 56 29
rect 60 19 64 29
rect 68 19 78 29
rect 92 19 96 29
rect 100 19 104 29
<< pdcontact >>
rect -17 72 -13 92
rect -9 72 -5 92
rect 4 72 8 92
rect 12 72 16 92
rect 20 72 24 92
rect 28 72 32 92
rect 36 72 40 92
rect 44 72 48 92
rect 52 72 56 92
rect 60 72 64 92
rect 68 72 78 92
rect 92 72 96 92
rect 100 72 104 92
<< psubstratepcontact >>
rect -17 8 104 14
<< nsubstratencontact >>
rect -17 97 104 103
<< polysilicon >>
rect -12 92 -10 94
rect -4 92 -2 94
rect 1 92 3 94
rect 9 92 11 94
rect 17 92 19 94
rect 25 92 27 94
rect 41 92 43 94
rect 49 92 51 94
rect 57 92 59 94
rect 65 92 67 94
rect 79 92 81 94
rect 84 92 86 94
rect 89 92 91 94
rect 97 92 99 94
rect -12 69 -10 72
rect -4 70 -2 72
rect -14 67 -10 69
rect -6 68 -2 70
rect -14 53 -12 67
rect -6 63 -4 68
rect -14 51 -10 53
rect -12 42 -10 51
rect -12 29 -10 38
rect -6 39 -4 59
rect 1 56 3 72
rect -6 37 -2 39
rect -4 29 -2 37
rect 1 29 3 52
rect 9 49 11 72
rect 17 63 19 72
rect 9 29 11 45
rect 17 29 19 59
rect 25 56 27 72
rect 41 63 43 72
rect 25 29 27 52
rect 41 29 43 59
rect 49 56 51 72
rect 49 29 51 52
rect 57 49 59 72
rect 57 29 59 45
rect 65 42 67 72
rect 79 68 81 72
rect 75 66 81 68
rect 75 49 77 66
rect 84 62 86 72
rect 82 60 86 62
rect 82 56 84 60
rect 89 56 91 72
rect 82 48 84 52
rect 82 46 86 48
rect 75 43 77 45
rect 75 41 81 43
rect 65 29 67 38
rect 79 29 81 41
rect 84 29 86 46
rect 89 29 91 52
rect 97 42 99 72
rect 97 29 99 38
rect -12 17 -10 19
rect -4 17 -2 19
rect 1 17 3 19
rect 9 17 11 19
rect 17 17 19 19
rect 25 17 27 19
rect 41 17 43 19
rect 49 17 51 19
rect 57 17 59 19
rect 65 17 67 19
rect 79 17 81 19
rect 84 17 86 19
rect 89 17 91 19
rect 97 17 99 19
<< polycontact >>
rect -8 59 -4 63
rect -14 38 -10 42
rect 0 52 4 56
rect 15 59 19 63
rect 8 45 12 49
rect 39 59 43 63
rect 25 52 29 56
rect 47 52 51 56
rect 55 45 59 49
rect 81 52 85 56
rect 89 52 93 56
rect 73 45 77 49
rect 63 38 67 42
rect 97 38 101 42
<< metal1 >>
rect -21 103 108 104
rect -21 97 -17 103
rect 104 97 108 103
rect -21 96 108 97
rect -9 92 -5 96
rect 20 92 24 96
rect 36 92 40 96
rect 52 92 56 96
rect 92 92 96 96
rect 12 69 16 72
rect 28 69 32 72
rect 12 66 32 69
rect 44 69 48 72
rect 60 69 64 72
rect 44 66 64 69
rect -4 59 15 63
rect 19 59 39 63
rect 43 59 93 63
rect 89 56 93 59
rect 4 52 25 56
rect 29 52 47 56
rect 51 52 81 56
rect 100 52 108 56
rect 100 49 104 52
rect 12 45 55 49
rect 59 45 73 49
rect 77 45 104 49
rect -10 38 4 42
rect 8 38 63 42
rect 76 38 97 42
rect 12 32 32 35
rect 12 29 16 32
rect 28 29 32 32
rect 44 32 64 35
rect 44 29 48 32
rect 60 29 64 32
rect -9 15 -5 19
rect 20 15 24 19
rect 36 15 40 19
rect 52 15 56 19
rect 92 15 96 19
rect -21 14 108 15
rect -21 8 -17 14
rect 104 8 108 14
rect -21 7 108 8
<< m2contact >>
rect -17 68 -13 72
rect 4 68 8 72
rect 68 68 78 72
rect 100 68 104 72
rect -21 52 -17 56
rect 4 38 8 42
rect 72 38 76 42
rect -17 29 -13 33
rect 4 29 8 33
rect 68 29 78 33
rect 100 29 104 33
<< metal2 >>
rect -17 33 -13 68
rect 4 42 8 68
rect 4 33 8 38
rect 68 33 72 68
rect 96 29 100 72
<< labels >>
rlabel nsubstratencontact 42 100 42 100 0 VDD
rlabel m2contact 102 31 102 31 0 S
rlabel metal2 -15 54 -15 54 0 Co
rlabel metal1 38 54 38 54 0 B
rlabel metal1 31 61 31 61 0 A
rlabel metal1 106 54 106 54 0 Ci
rlabel psubstratepcontact 43 10 43 10 0 GND
<< end >>
