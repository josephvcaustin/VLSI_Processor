magic
tech scmos
timestamp 1481316034
<< metal1 >>
rect 0 94 87 95
rect 28 89 30 91
rect -3 49 4 53
rect 80 49 83 55
rect -3 42 8 46
rect 28 9 30 11
rect 0 5 87 6
<< m2contact >>
rect -3 57 1 61
rect 32 49 36 53
rect 68 49 72 53
rect 32 42 36 46
rect 60 42 64 46
rect -3 34 1 38
rect 24 25 28 29
rect 52 17 56 21
<< metal2 >>
rect 1 57 36 61
rect 32 53 36 57
rect 32 38 36 42
rect 1 34 36 38
rect 60 29 64 42
rect 28 25 64 29
rect 68 21 72 49
rect 56 17 72 21
use nand  nand_0
timestamp 1480790700
transform 1 0 23 0 1 67
box -23 -61 8 27
use nand  nand_1
timestamp 1480790700
transform 1 0 51 0 1 67
box -23 -61 8 27
use nand  nand_2
timestamp 1480790700
transform 1 0 79 0 1 67
box -23 -61 8 27
<< labels >>
rlabel m2contact -1 59 -1 59 1 D
rlabel m2contact -1 36 -1 36 1 Clk
rlabel metal1 -1 51 -1 51 1 A
rlabel metal1 -1 44 -1 44 1 Clk_
rlabel metal1 28 89 30 91 1 VDD
rlabel metal1 28 9 30 11 1 GND
rlabel metal1 81 53 81 53 1 En
<< end >>
